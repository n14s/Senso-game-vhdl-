library ieee; use ieee.std_logic_1164.all;
entity input is
end entity input;
