entity tb is
--TB entity bleibt leer
end entity tb;