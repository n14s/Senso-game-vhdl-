library ieee; use ieee.std_logic_1154.all;
