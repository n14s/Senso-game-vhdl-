root@nikx.4606:1574890555