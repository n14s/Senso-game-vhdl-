library ieee; use ieee.std_logic_1164.all;

architecture behav of input is
begin
end architecture behav;